library ieee;
use ieee.std_logic.1164.all
